`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    21:08:04 11/17/2016 
// Design Name: 
// Module Name:    ALU16 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module ALU16(
    input [16:0] x,
    input [16:0] y,
    output [16:0] out,
    input cin,
    output cout,
    output lt,
    output eq,
    output gt,
    output v,
    input [2:0] opcode
    );


endmodule
